// Top level file for USB RX
